localparam  int OBJECT_WIDTH_X = 50;
localparam  int OBJECT_HEIGHT_Y = 50;

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h69, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h64, 8'h68, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h8D, 8'hB2, 8'hB1, 8'h8D, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h8D, 8'hB1, 8'h8D, 8'h68, 8'h64, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h91, 8'h64, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h64, 8'h64, 8'h64, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'h8D, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'hC8, 8'hC8, 8'hC8, 8'hC8, 8'hCD, 8'hCD, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hCD, 8'hC9, 8'hC8, 8'hC8, 8'h88, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h8C, 8'h8C, 8'h68, 8'h84, 8'h84, 8'hA4, 8'hA4, 8'hC4, 8'hC4, 8'hC8, 8'hE8, 8'hCD, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hE8, 8'hE8, 8'hC4, 8'hA4, 8'h84, 8'h88, 8'h8C, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h8C, 8'h90, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h64, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h84, 8'hA4, 8'hC8, 8'hC4, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'hE8, 8'h84, 8'h80, 8'h80, 8'h88, 8'hF8, 8'hF8, 8'h44, 8'h90, 8'hD4, 8'hD4, 8'hF8, 8'h6C, 8'h24, 8'hF8, 8'hF8, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h64, 8'h80, 8'h80, 8'h80, 8'h80, 8'hA4, 8'hC8, 8'hC8, 8'hC8, 8'hE8, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'hC8, 8'h80, 8'h80, 8'h68, 8'hD4, 8'hFC, 8'hB0, 8'hD8, 8'hD4, 8'hD8, 8'hF8, 8'hB4, 8'h90, 8'hF8, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hC8, 8'hC4, 8'hC4, 8'hA4, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE8, 8'hC4, 8'h60, 8'h68, 8'h8C, 8'hB0, 8'hD4, 8'hB0, 8'h8C, 8'h8C, 8'h8C, 8'hB0, 8'hB0, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h8C, 8'h64, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hA4, 8'h80, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hC8, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h84, 8'h80, 8'h84, 8'hC8, 8'h84, 8'h80, 8'h80, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h88, 8'h6C, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h60, 8'hC4, 8'hC4, 8'h80, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h6C, 8'h88, 8'hC8, 8'h84, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h88, 8'hC8, 8'h84, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h8C, 8'h8C, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h68, 8'hA8, 8'hA4, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h90, 8'h90, 8'h90, 8'hB4, 8'hB5, 8'hD9, 8'hFD, 8'hFD, 8'h90, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h6C, 8'h88, 8'hA8, 8'hA4, 8'h60, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h68, 8'h68, 8'h68, 8'h68, 8'hB0, 8'hD9, 8'hB5, 8'hD9, 8'hD5, 8'h8C, 8'hB5, 8'hB4, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h88, 8'hA8, 8'h84, 8'h60, 8'h80, 8'h89, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h88, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h48, 8'h25, 8'h29, 8'h49, 8'h84, 8'h80, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h8C, 8'h88, 8'h68, 8'h24, 8'h29, 8'h25, 8'h29, 8'h49, 8'hA8, 8'hA4, 8'h84, 8'h80, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h88, 8'h8C, 8'h8C, 8'h8C, 8'h88, 8'h68, 8'h68, 8'h44, 8'h24, 8'h24, 8'h48, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hC8, 8'hA4, 8'h80, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8C, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h48, 8'h48, 8'h44, 8'h44, 8'h48, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'hC8, 8'hA4, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hC8, 8'hA4, 8'h80, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h69, 8'h8D, 8'h6D, 8'h6D, 8'h8D, 8'h8D, 8'h6C, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hE8, 8'h84, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h49, 8'h72, 8'h72, 8'h4E, 8'h9A, 8'h91, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hC8, 8'hA4, 8'h80, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6D, 8'h6D, 8'h4E, 8'h72, 8'h72, 8'h76, 8'h96, 8'h96, 8'h96, 8'h9A, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hA8, 8'hE8, 8'h84, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h6E, 8'h92, 8'h93, 8'h76, 8'h76, 8'h96, 8'hBF, 8'hBF, 8'hBF, 8'h9A, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h88, 8'hE8, 8'hA4, 8'h60, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h4D, 8'h6D, 8'h8D, 8'h92, 8'h93, 8'h93, 8'h93, 8'h72, 8'h77, 8'h76, 8'h76, 8'h76, 8'h72, 8'h6D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hE8, 8'hC4, 8'h80, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h4E, 8'h6D, 8'h89, 8'h6D, 8'h92, 8'h92, 8'h8E, 8'h72, 8'h72, 8'h72, 8'h71, 8'h6D, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'hC8, 8'hC8, 8'h80, 8'h89, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h64, 8'hA4, 8'hC8, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h91, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h6C, 8'h6C, 8'h6C, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h80, 8'hA4, 8'hE8, 8'h84, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h88, 8'h88, 8'h8C, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h64, 8'h80, 8'h84, 8'hE8, 8'h84, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB1, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hFF, 8'hFF, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h84, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hA4, 8'h80, 8'h89, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h6C, 8'h68, 8'h8D, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h64, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hA4, 8'h80, 8'h84, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h8D, 8'h91, 8'h91, 8'h6C, 8'h68, 8'h6C, 8'hFF, 8'hFF, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h8C, 8'h68, 8'h68, 8'h6C, 8'h64, 8'h80, 8'h80, 8'h80, 8'h80, 8'hA4, 8'hC4, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'hA4, 8'hC8, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h84, 8'hC8, 8'h80, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h64, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h84, 8'hC8, 8'h84, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h68, 8'h68, 8'h88, 8'h88, 8'h88, 8'h88, 8'h68, 8'h68, 8'h68, 8'h64, 8'h64, 8'h64, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'h84, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h91, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h84, 8'h80, 8'h80, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h6C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'h84, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h68, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h84, 8'h80, 8'h80, 8'h68, 8'h8C, 8'h68, 8'h88, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h68, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hA4, 8'h80, 8'hB2, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h84, 8'h84, 8'h84, 8'h68, 8'h6C, 8'h88, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h84, 8'h84, 8'h84, 8'h80, 8'h80, 8'h80, 8'h80, 8'hC8, 8'hC4, 8'h60, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hA8, 8'hE8, 8'hE8, 8'h88, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hC8, 8'hE8, 8'hE8, 8'hC8, 8'hC4, 8'hA4, 8'hA4, 8'hC8, 8'hC8, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'hD1, 8'hD1, 8'h8D, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hAD, 8'hD1, 8'hCD, 8'hCD, 8'hC8, 8'hE8, 8'hC8, 8'hC8, 8'hE8, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h88, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h91, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hC8, 8'hE8, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'hFF, 8'hFF, 8'h8D, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h68, 8'h8C, 8'h8D, 8'hB1, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h8C, 8'h91, 8'hFF, 8'hFF, 8'hB1, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8C, 8'h8C, 8'h8D, 8'h91, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h6C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'h68, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h68, 8'h68, 8'h8C, 8'h91, 8'hFF, 8'hFF, 8'h8D, 8'h68, 8'h68, 8'h68, 8'h8D, 8'h91, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h91, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};

wire [7:0] red_sig, green_sig, blue_sig;
assign red_sig     = {object_colors[offsetY][offsetX][7:5] , 5'd0};
assign green_sig   = {object_colors[offsetY][offsetX][4:2] , 5'd0};
assign blue_sig    = {object_colors[offsetY][offsetX][1:0] , 6'd0};


