module NumbersBitMap	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] offsetX,// offset from top left  position 
					input 	logic	[10:0] offsetY,
					input		logic	InsideRectangle, //input that the pixel is within a bracket 
					input 	logic	[9:0] score, // digits to display
					input		logic [1:0] lives  ,
					
					output	logic				drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0]		RGBout
);
// generating a smily bitmap 

parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 
localparam  int LIFE_WIDTH_X = 32;
localparam  int LIFE_HEIGHT_Y = 32;
localparam  int SCORE_WIDTH_X = 32;
localparam  int SCORE_HEIGHT_Y = 96;
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 					

int digits[2:0] ;
int num ;


bit [0:15] [0:31] [0:15] number_bitmap  = {


{16'b	0000001111100000,
16'b	0000111111111000,
16'b	0000111111111000,
16'b	0001111111111100,
16'b	0011111001111100,
16'b	0011100000111110,
16'b	0111100000011110,
16'b	0111100000011110,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000011110,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111110000111100,
16'b	0011111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111110000,
16'b	0000011111000000},
																	
{16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000011111100000,
16'b	0000111111100000,
16'b	0001111111100000,
16'b	0011111111100000,
16'b	0111111011100000,
16'b	0111100011100000,
16'b	0111000011100000,
16'b	0010000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111},
																	
{16'b	0000111111100000,
16'b	0001111111110000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000011111100,
16'b	1110000001111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0011111000000000,
16'b	0111110000000001,
16'b	1111100000000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},
																	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000001111100,
16'b	1110000001111100,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0001111111110000,
16'b	0001111111000000,
16'b	0001111111111000,
16'b	0001111111111000,
16'b	0000000011111100,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000111111,
16'b	1110000001111110,
16'b	1111100011111110,
16'b	1111111111111100,
16'b	1111111111111000,
16'b	0111111111111000,
16'b	0001111111000000},
																	
{16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000111111000,
16'b	0000001111111000,
16'b	0000001101111000,
16'b	0000011101111000,
16'b	0000011101111000,
16'b	0000111101111000,
16'b	0001111101111000,
16'b	0001111101111000,
16'b	0001111001111000,
16'b	0011111001111000,
16'b	0011110001111000,
16'b	0111100001111000,
16'b	0111100001111000,
16'b	1111000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000011111100},
																	
{16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111110,
16'b	0111111111111100,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111111111100000,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0010000011111110,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	1000000000111110,
16'b	1100000001111110,
16'b	1111100011111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	0001111111000000},
																	
{16'b	0000000111111100,
16'b	0000011111111110,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0001111100001111,
16'b	0011111100000001,
16'b	0011111000000000,
16'b	0111110000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111001111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	1111111111111111,
16'b	1111111101111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111100000001111,
16'b	1111100000001111,
16'b	0111110000011111,
16'b	0111111101111110,
16'b	0011111111111110,
16'b	0001111111111100,
16'b	0001111111111000,
16'b	0000011111100000},
																	
{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1100000000001111,
16'b	1000000000011111,
16'b	0000000000011111,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000000111100000,
16'b	0000001111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000011110000000,
16'b	0000111110000000,
16'b	0000111100000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0001111100000000},
																	
{16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111111111110,
16'b	0111111011111110,
16'b	1111100000111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111100000,
16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111001111110,
16'b	1111100000111111,
16'b	1111000000001111,
16'b	1110000000001111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111001111111,
16'b	1111111111111110,
16'b	0111111111111110,
16'b	0011111111111000,
16'b	0001111111110000},
																	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0011111111111000,
16'b	0111111111111100,
16'b	1111111011111100,
16'b	1111100000111110,
16'b	1111000000011110,
16'b	1111000000011111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111011111111,
16'b	1111111111111111,
16'b	0111111111111111,
16'b	0011111111111111,
16'b	0001111111001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011110,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000001111100,
16'b	1000000011111100,
16'b	1111000011111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111100000,
16'b	0011111100000000},

{16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000111111110000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0001110000111100,
16'b	0001100000011100,
16'b	0011100000011100,
16'b	0011000000001100,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111},


{16'b	1111111111110000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	0111000011111110,
16'b	0111000000111111,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000001111100,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111100000,
16'b	0111111111110000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0111000001111110,
16'b	0111000000111111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000000111,
16'b	0111000000000111,
16'b	0111000000001111,
16'b	0111000000011111,
16'b	0111000001111111,
16'b	1111111111111110,
16'b	1111111111111110,
16'b	1111111111111000,
16'b	1111111111110000},

{16'b	0000001111111000,
16'b	0000111111111100,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0011111001000011,
16'b	0011100000000001,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111100000000000,
16'b	0111110000000000,
16'b	0111110000000001,
16'b	0011111001000011,
16'b	0011111111111111,
16'b	0001111111111110,
16'b	0000111111111100,
16'b	0000011111111000},


{16'b	1111111111100000,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	0111000001111100,
16'b	0111000000111110,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000000111100,
16'b	0111000001111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111000000},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000001000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000}



} ;
logic [0:LIFE_HEIGHT_Y-1] [0:LIFE_WIDTH_X-1] [8-1:0] life_colors = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h45, 8'h6D, 8'hB6, 8'h68, 8'h20, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h44, 8'h04, 8'h68, 8'hA8, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h88, 8'h44, 8'h44, 8'hCC, 8'h64, 8'h6D, 8'hFF, 8'hBA, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'hCC, 8'h68, 8'hCC, 8'hCC, 8'h24, 8'h25, 8'h49, 8'h44, 8'h64, 8'h44, 8'h49, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hA8, 8'h44, 8'h92, 8'hBA, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h25, 8'hA8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h44, 8'h44, 8'h44, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hAC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h44, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h04, 8'h05, 8'h24, 8'hAC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hAC, 8'hA8, 8'h8C, 8'hAD, 8'hAD, 8'h88, 8'hAC, 8'hCC, 8'hCC, 8'hCC, 8'hAC, 8'h64, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h09, 8'h0E, 8'h04, 8'hA8, 8'hCC, 8'hCC, 8'hAC, 8'h88, 8'hAD, 8'hD1, 8'hF6, 8'hF6, 8'hF6, 8'h8D, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h20, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h09, 8'h0E, 8'h12, 8'h09, 8'h24, 8'h44, 8'h68, 8'hB1, 8'hD5, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hAD, 8'h88, 8'hA8, 8'hCC, 8'hCC, 8'hCC, 8'h44, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h09, 8'h0E, 8'h32, 8'h32, 8'h0E, 8'h00, 8'hB1, 8'hF6, 8'hF6, 8'hF5, 8'hD5, 8'hF5, 8'hF6, 8'hAD, 8'hB1, 8'h89, 8'hCC, 8'hCC, 8'hCC, 8'hA8, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h04, 8'h09, 8'h09, 8'h0E, 8'h32, 8'h12, 8'h49, 8'hB2, 8'hB1, 8'hD1, 8'hB1, 8'hB6, 8'hB2, 8'hD1, 8'hF6, 8'hD1, 8'hAC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h20, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h92, 8'h04, 8'h09, 8'h09, 8'h05, 8'h09, 8'h29, 8'hDB, 8'hFF, 8'hDB, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hD5, 8'hAD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h24, 8'h05, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h6D, 8'h05, 8'h09, 8'h05, 8'h09, 8'h05, 8'h6D, 8'hFF, 8'hDB, 8'hFF, 8'hB6, 8'hFF, 8'hDA, 8'hFF, 8'hDB, 8'hB1, 8'hAC, 8'hAC, 8'hAC, 8'hCC, 8'hCC, 8'hAC, 8'h04, 8'h09, 8'h05, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h6D, 8'h09, 8'h0E, 8'h0E, 8'h09, 8'h05, 8'h49, 8'hDB, 8'hDB, 8'h91, 8'h91, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hD1, 8'h68, 8'hAD, 8'h8D, 8'hAC, 8'hCC, 8'h44, 8'h05, 8'h0E, 8'h09, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h6D, 8'h09, 8'h0E, 8'h12, 8'h32, 8'h32, 8'h09, 8'h8D, 8'hB1, 8'hD5, 8'hD1, 8'hB2, 8'hDA, 8'hB6, 8'hB1, 8'hF5, 8'hB1, 8'hB1, 8'hB1, 8'h89, 8'h44, 8'h00, 8'h09, 8'h09, 8'h09, 8'h04, 8'h24, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h6D, 8'h04, 8'h0E, 8'h0E, 8'h0E, 8'h32, 8'h29, 8'hB1, 8'hD5, 8'hD5, 8'hF6, 8'hF5, 8'hD1, 8'hD1, 8'hF6, 8'hF6, 8'hF6, 8'hD5, 8'h8D, 8'h00, 8'h04, 8'h09, 8'h09, 8'h09, 8'h09, 8'h05, 8'h00, 8'hDB, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h05, 8'h09, 8'h09, 8'h09, 8'h05, 8'h8D, 8'hB1, 8'hD1, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF5, 8'h44, 8'h04, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h05, 8'h00, 8'hB6, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h05, 8'h09, 8'h09, 8'h05, 8'h69, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hD1, 8'h00, 8'h36, 8'h37, 8'h36, 8'h32, 8'h0E, 8'h0E, 8'h0D, 8'h09, 8'h00, 8'h92, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h09, 8'h09, 8'h49, 8'hF5, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hD1, 8'h00, 8'h09, 8'h2E, 8'h32, 8'h32, 8'h32, 8'h12, 8'h0E, 8'h0E, 8'h05, 8'h92, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h09, 8'h09, 8'h69, 8'hD1, 8'hD5, 8'hD5, 8'hD1, 8'hD1, 8'hB1, 8'hB1, 8'hB1, 8'hF6, 8'hF6, 8'hB1, 8'h00, 8'h04, 8'h05, 8'h05, 8'h09, 8'h09, 8'h0E, 8'h0E, 8'h0E, 8'h05, 8'h92, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h04, 8'h09, 8'h05, 8'h04, 8'h24, 8'h25, 8'h24, 8'h8D, 8'hD1, 8'hD5, 8'hF5, 8'hF6, 8'hF6, 8'hB1, 8'h40, 8'h00, 8'h05, 8'h09, 8'h05, 8'h05, 8'h09, 8'h09, 8'h09, 8'h04, 8'hB6, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h05, 8'h09, 8'h09, 8'h09, 8'h12, 8'h05, 8'h20, 8'hD1, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hB1, 8'h84, 8'h60, 8'h00, 8'h2E, 8'h09, 8'h09, 8'h09, 8'h09, 8'h05, 8'h04, 8'hDB, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h05, 8'h09, 8'h0E, 8'h05, 8'h20, 8'h84, 8'hAD, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hB1, 8'h64, 8'h84, 8'h20, 8'h00, 8'h09, 8'h0E, 8'h09, 8'h09, 8'h05, 8'h49, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h09, 8'h05, 8'h00, 8'h64, 8'h84, 8'h8D, 8'hB1, 8'hD1, 8'hD1, 8'hB1, 8'h91, 8'h64, 8'h84, 8'h64, 8'h60, 8'h00, 8'h05, 8'h0E, 8'h09, 8'h04, 8'hB6, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h00, 8'h64, 8'h84, 8'h84, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hDB, 8'h84, 8'h84, 8'h64, 8'h84, 8'h84, 8'h20, 8'h05, 8'h09, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h40, 8'h84, 8'h84, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h84, 8'h84, 8'h64, 8'h84, 8'h84, 8'h84, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h20, 8'h44, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h84, 8'h84, 8'h64, 8'h84, 8'h84, 8'h40, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h49, 8'h00, 8'h24, 8'h6D, 8'h92, 8'hB6, 8'hDA, 8'h92, 8'h64, 8'h84, 8'h40, 8'h20, 8'h00, 8'h49, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'h92, 8'h92, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};
logic [0:SCORE_HEIGHT_Y-1] [0:SCORE_WIDTH_X-1] [8-1:0] score_colors = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h49, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h49, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h49, 8'hB6, 8'hDA, 8'hDA, 8'hB6, 8'h6D, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h24, 8'hDA, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h49, 8'h00, 8'h00, 8'h24, 8'hDB, 8'h49, 8'h00, 8'h00, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h24, 8'h24, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'h92, 8'h24, 8'h00, 8'h24, 8'h92, 8'hFF, 8'hDB, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'h92, 8'h92, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h49, 8'h00, 8'h24, 8'h00, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'h92, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'hDA, 8'hFF, 8'h92, 8'h00, 8'h25, 8'h92, 8'h49, 8'h00, 8'hB6, 8'hFF, 8'h49, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'h92, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h24, 8'hFF, 8'hFF, 8'h24, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h6D, 8'h123, 8'h92, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h24, 8'h00, 8'h00, 8'h25, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h24, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h24, 8'h00, 8'h00, 8'h00, 8'h25, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h24, 8'hFF, 8'hDB, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'hB6, 8'hFF, 8'h92, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h24, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h92, 8'h25, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'h6D, 8'hDB, 8'h49, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h24, 8'hFF, 8'hDB, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'h6D, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'hDA, 8'hFF, 8'h25, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h6D, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h6D, 8'h123, 8'hB6, 8'h00, 8'h24, 8'h92, 8'hDA, 8'hDA, 8'h92, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h92, 8'hFF, 8'hDB, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h6D, 8'h00, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hB6, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hDB, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h24, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h00, 8'h49, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h92, 8'hFF, 8'h24, 8'h00, 8'h49, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hDB, 8'hB6, 8'h49, 8'h24, 8'h00, 8'h25, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'hB6, 8'hFF, 8'hDB, 8'h92, 8'h6D, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6D, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'hB6, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h92, 8'hDA, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h24, 8'h24, 8'h00, 8'h24, 8'h49, 8'h92, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h6D, 8'hFF, 8'h123, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h92, 8'hDB, 8'h24, 8'h00, 8'h49, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h49, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hDA, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h24, 8'h00, 8'h6D, 8'h123, 8'h92, 8'h00, 8'h00, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'h92, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h6D, 8'hDB, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h49, 8'hFF, 8'hB6, 8'h6D, 8'hDB, 8'hFF, 8'h24, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'h6D, 8'h24, 8'h00, 8'h25, 8'h6D, 8'hB6, 8'h25, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h24, 8'h24, 8'h49, 8'h92, 8'hB6, 8'h92, 8'h25, 8'h00, 8'h24, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hDA, 8'h24, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h49, 8'h92, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h49, 8'h24, 8'h00, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'hB6, 8'h123, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h49, 8'h00, 8'h00, 8'h25, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h24, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'hDB, 8'hDB, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h92, 8'hFF, 8'h6D, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hDA, 8'hDA, 8'hDA, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h92, 8'h92, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h24, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h24, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h24, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h24, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h49, 8'h49, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'h24, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h92, 8'h123, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h25, 8'h00, 8'h00, 8'h49, 8'h00, 8'h24, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h6D, 8'hFF, 8'h49, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h24, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'hB6, 8'hFF, 8'h25, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hB6, 8'hDB, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'hDB, 8'h49, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h24, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hB6, 8'h24, 8'h00, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h49, 8'h24, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};
// pipeline (ff) to get the pixel color from the array 	 
	
// LifeBitMap														   
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		drawingRequest <=	1'b0;
	end
	else begin
	if (offsetX<96) begin //life , score , numbers
	for (int i=0;i<lives;i++) begin
		if (InsideRectangle == 1'b1)  // inside an external bracket 
			RGBout <= life_colors[offsetY][offsetX+i*32];	//get RGB from the colors table  0 - 
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
		end
		end
	else if(offsetX<192) begin
		if (InsideRectangle == 1'b1)  // inside an external bracket 
			RGBout <= score_colors[offsetY][offsetX+192];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end
	else begin
		num <= score ;
	
	for (int i=0;i<3;i++)
	begin
			digits[i] <= num % 10 ;
			drawingRequest <= (number_bitmap[digits[2-i]][offsetY][offsetX+192+i*32]) && (InsideRectangle == 1'b1 );
			RGBout <= digit_color ;
			num <= num / 10 ;
	end
	end 
	end
	end	// ScoreBitMap														   
/*always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1)  // inside an external bracket 
			RGBout <= score_colors[offsetY][offsetX];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
		end
		end
	end 
end	*/
														
												


// NumbersBitMap
/*always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
	end
	else begin
	for (int i=0;i<3;i++)
	{
			drawingRequest <= (number_bitmap[score[i][3:0]][offsetY][offsetX<<i]) && (InsideRectangle == 1'b1 );
	}
	end 
end

assign RGBout = digit_color ; // this is a fixed color
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap
*/
endmodule