module	controller (	
					input logic clk ,
					input logic resetN 
);

always_ff@(posedge clk or negedge resetN)
begin
	//if(!resetN)	
		
	//else 
	//begin 
	
		
	//end
end 
endmodule 