module	StartBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket
					
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
);	
// generating a bolt bitmap 						

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 						 
localparam  int OBJECT_WIDTH_X = 64;
localparam  int OBJECT_HEIGHT_Y = 64;

logic [0:OBJECT_HEIGHT_Y-1] [1*64-1:0] object_colors = {
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000111100000000000000000000111100000000000000000},
{64'b0000000000000000000111100000000000000000000111100000000000000000},
{64'b0000000000000000000111100000000000000000000111100000000000000000},
{64'b0000000000000000000111100000000000000000000111100000000000000000},
{64'b0000000000000000000000011110000000000001111000000000000000000000},
{64'b0000000000000000000000011110000000000001111000000000000000000000},
{64'b0000000000000000000000011110000000000001111000000000000000000000},
{64'b0000000000000000000000011110000000000001111000000000000000000000},
{64'b0000000000000000000111111111111111111111111111100000000000000000},
{64'b0000000000000000000111111111111111111111111111100000000000000000},
{64'b0000000000000000000111111111111111111111111111100000000000000000},
{64'b0000000000000000000111111111111111111111111111100000000000000000},
{64'b0000000000000001111111100001111111111110000111111110000000000000},
{64'b0000000000000001111111100001111111111110000111111110000000000000},
{64'b0000000000000001111111100001111111111110000111111110000000000000},
{64'b0000000000000001111111100001111111111110000111111110000000000000},
{64'b0000000000011111111111111111111111111111111111111111111000000000},
{64'b0000000000001111111111111111111111111111111111111111111000000000},
{64'b0000000000011111111111111111111111111111111111111111111000000000},
{64'b0000000000011111111111111111111111111111111111111111111000000000},
{64'b0000000000011110000111111111111111111111111111100001111000000000},
{64'b0000000000011110000111111111111111111111111111100001111000000000},
{64'b0000000000011110000111111111111111111111111111100001111000000000},
{64'b0000000000011110000111111111111111111111111111100001111000000000},
{64'b0000000000011110000111100000000000000000000111100001111000000000},
{64'b0000000000011110000111100000000000000000000111100001111000000000},
{64'b0000000000011110000111100000000000000000000111100001111000000000},
{64'b0000000000001110000011100000000000000000000111100001110000000000},
{64'b0000000000000000000000011111111000011111111000000000000000000000},
{64'b0000000000000000000000011111111000011111111000000000000000000000},
{64'b0000000000000000000000011111111000011111111000000000000000000000},
{64'b0000000000000000000000001111111000001110010000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0011111001111001111100111000110000001110011110001100011110011111},
{64'b0011001101000101100001001101001000010010001100001100010001000100},
{64'b0011001101100101100001100001000000011000001100010110010011000100},
{64'b0011000001101101100000011000011000000110001100011110011011000100},
{64'b0011000001000101100001001101001000010011001100110010010001000100},
{64'b0011000001000101111100111001111000011110001000110011010001000100},
{64'b0000000000000000000000000000000000000000000000000000000000000000},
{64'b0000000000000000000000000000000000000000000000000000000000000000}
};

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1)  // inside an external bracket 
			RGBout <= object_colors[offsetY][offsetX];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule

