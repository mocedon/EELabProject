module	EndBitBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket
					
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
);	
// generating a bolt bitmap 						

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 						 
localparam  int OBJECT_WIDTH_X = 32;
localparam  int OBJECT_HEIGHT_Y = 32;

logic [0:OBJECT_HEIGHT_Y-1] [1*32-1:0] object_colors = {
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000111100111001111110001110000},
{32'b00001111001111101111111011100000},
{32'b00001100001101101101011011000000},
{32'b00001101101111101101011011110000},
{32'b00001101101111101101011011000000},
{32'b00001111101101101101011011100000},
{32'b00000111001101101001001001110000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000111001101101111001111100000},
{32'b00001111101101101110011111110000},
{32'b00001101101101101100011000110000},
{32'b00001101101101101111011111110000},
{32'b00001101101111101100011111100000},
{32'b00001111100111001110011001110000},
{32'b00000111000010001111011000110000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b00000000000000000000000000000000},
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111},
{32'b11111111111111111111111111111111}
};
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1)  // inside an external bracket 
			RGBout <= object_colors[offsetY][offsetX];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule
